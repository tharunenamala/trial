module simple;
intial
begin
$display()
endmodule
